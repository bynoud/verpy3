
module modname();
endmodule
