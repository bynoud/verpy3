
module legacy_direct (); endmodule
